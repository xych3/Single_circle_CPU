`timescale 1ns / 1ps
module InsMem(
    input RW,                   // read or write
    input [7:0] IAddr,          // instruction address
    output reg [31:0] IDataOut  // instruction output
    );
    reg [7:0] Inst[0:255];      // Instructions(21) reg(8) - 21*4=84
    always @(IAddr) begin
        IDataOut = {Inst[IAddr],Inst[IAddr+1],Inst[IAddr+2],Inst[IAddr+3]};
    end

    initial begin
        {Inst[0],Inst[1],Inst[2],Inst[3]} <= 32'b000000001000_00000_000_00001_0010011;          // 0x0000_0000
        {Inst[4],Inst[5],Inst[6],Inst[7]} <= 32'b000000000010_00000_110_00010_0010011;          // 0x0000_0004
        {Inst[8],Inst[9],Inst[10],Inst[11]} <= 32'b0000000_00001_00010_000_00011_0110011;       // 0x0000_0008
        {Inst[12],Inst[13],Inst[14],Inst[15]} <= 32'b0100000_00010_00011_000_00101_0110011;     // 0x0000_000C
        {Inst[16],Inst[17],Inst[18],Inst[19]} <= 32'b0000000_00010_00101_111_00100_0110011;     // 0x0000_0010
        {Inst[20],Inst[21],Inst[22],Inst[23]} <= 32'b0000000_00010_00110_110_01000_0110011;     // 0x0000_0014
        {Inst[24],Inst[25],Inst[26],Inst[27]} <= 32'b000000000001_01000_001_01000_0010011;      // 0x0000_0018
        {Inst[28],Inst[29],Inst[30],Inst[31]} <= 32'b1_111111_00001_01000_001_1110_1_1100011;   // 0x0000_001C
        {Inst[32],Inst[33],Inst[34],Inst[35]} <= 32'b000000000100_00010_010_00110_0010011;      // 0x0000_0020
        {Inst[36],Inst[37],Inst[38],Inst[39]} <= 32'b000000000000_00110_010_00111_0010011;      // 0x0000_0024
        {Inst[40],Inst[41],Inst[42],Inst[43]} <= 32'b000000001000_00111_000_00111_0010011;      // 0x0000_0028
        {Inst[44],Inst[45],Inst[46],Inst[47]} <= 32'b1_111111_00001_00111_000_1110_1_1100011;   // 0x0000_002C
        {Inst[48],Inst[49],Inst[50],Inst[51]} <= 32'b0000000_00010_00001_010_00100_0100011;     // 0x0000_0030
        {Inst[52],Inst[53],Inst[54],Inst[55]} <= 32'b000000000100_00001_010_01001_0000011;      // 0x0000_0034
        {Inst[56],Inst[57],Inst[58],Inst[59]} <= 32'b111111111110_00000_000_01010_0010011;      // 0x0000_0038
        {Inst[60],Inst[61],Inst[62],Inst[63]} <= 32'b000000000001_01010_000_01010_0010011;      // 0x0000_003C
        {Inst[64],Inst[65],Inst[66],Inst[67]} <= 32'b1_111111_00000_01010_100_1110_1_1100011;   // 0x0000_0040
        {Inst[68],Inst[69],Inst[70],Inst[71]} <= 32'b000000000010_00010_111_01011_0010011;      // 0x0000_0044
        {Inst[72],Inst[73],Inst[74],Inst[75]} <= 32'b0_0000000100_0_00000000_01000_1101111;     // 0x0000_0048
        {Inst[76],Inst[77],Inst[78],Inst[79]} <= 32'b0000000_00010_00100_110_01000_0110011;     // 0x0000_004C
        {Inst[80],Inst[81],Inst[82],Inst[83]} <= 32'b000000000000_xxxxx_000_xxxxx_1110011;      // 0x0000_0050
    end
endmodule
